`include "uart_top_monitor.sv"
`include "uart_top_driver.sv"
`include "uart_top_sequencer.sv"
`include "uart_top_agent.sv"