`include "uart_monitor.sv"
`include "uart_driver.sv"
`include "uart_sequencer.sv"
`include "uart_agent.sv"